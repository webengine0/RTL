`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    10:29:11 10/15/2024 
// Design Name: 
// Module Name:    PC_Adder 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module PC_Adder(a,b,c
    );
	 input [31:0]a,b;
	 output [31:0]c;
	 
	 assign c = a + b; 


endmodule
